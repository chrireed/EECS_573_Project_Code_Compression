//TODO: Make the logic here combinational (for a preloaded dictionary, we don't need this to be clocked...)
//We can make use of that saved cycle though.

//Inputs:
//key_data_in: Compressed key (index into LUT)
//val_lookup_in: Enter an uncompressed bitstring, returns existence in val_lookup_res.
module dictionary #(
  parameter KEY_WIDTH  = 4,
  parameter VAL_WIDTH  = 8)
  (
  //------------Input Ports--------------                        
  input  [KEY_WIDTH-1:0]   key_lookup_in, //Lookup this key (index bits / compressed bits)
  input  [VAL_WIDTH-1:0]   val_lookup_in, //lookup this value (uncompressed bits for field)
  //----------Output Ports--------------
  output reg [VAL_WIDTH-1:0]   val_out,  // found this value (uncompressed bits) for the compressed bits given.
  output reg [KEY_WIDTH-1:0]   key_out,  // found this value (compressed bits) for the uncompressed bits given.
  output reg                   val_lookup_result  //is the uncompressed bits an entry in the table?
  //------------Internal Variables--------
  );
  // Stored CAM memory (KEY_WIDTH entries, each 8-bit wide)
  reg [VAL_WIDTH-1:0] memory [2**KEY_WIDTH - 1:0];

  integer i;

  initial begin
    val_lookup_result = 1'b0;
    val_out <= {VAL_WIDTH{1'b0}};  // VAL_WIDTH-bit zero

    //insert mem init stuff here
    for (i = 0; i < 2**KEY_WIDTH; i = i + 1) begin
      memory[i] = i + 1; // Each memory location is filled with its index value
    end
  end

  always @* begin
      val_out = memory[key_lookup_in];
      val_lookup_result = 1'b0;  
      key_out = 0;                  
      
      for (i = 0; i < (2**KEY_WIDTH); i = i + 1) begin
          if (memory[i] == val_lookup_in && ~val_lookup_result) begin
              val_lookup_result = 1'b1;
              key_out = i;   
          end
      end
  end

endmodule